VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cla
  CLASS BLOCK ;
  FOREIGN cla ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 32.680 500.000 33.280 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 94.560 500.000 95.160 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 156.440 500.000 157.040 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 218.320 500.000 218.920 ;
    END
  END A[3]
  PIN B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 280.200 500.000 280.800 ;
    END
  END B[0]
  PIN B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 342.080 500.000 342.680 ;
    END
  END B[1]
  PIN B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 403.960 500.000 404.560 ;
    END
  END B[2]
  PIN B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 465.840 500.000 466.440 ;
    END
  END B[3]
  PIN S[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END S[0]
  PIN S[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END S[3]
  PIN cin
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END cin
  PIN cout
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END cout
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 5.520 10.640 494.040 487.120 ;
      LAYER met2 ;
        RECT 7.910 10.695 492.560 487.065 ;
      LAYER met3 ;
        RECT 4.000 466.840 496.000 487.045 ;
        RECT 4.000 465.440 495.600 466.840 ;
        RECT 4.000 458.000 496.000 465.440 ;
        RECT 4.400 456.600 496.000 458.000 ;
        RECT 4.000 404.960 496.000 456.600 ;
        RECT 4.000 403.560 495.600 404.960 ;
        RECT 4.000 375.040 496.000 403.560 ;
        RECT 4.400 373.640 496.000 375.040 ;
        RECT 4.000 343.080 496.000 373.640 ;
        RECT 4.000 341.680 495.600 343.080 ;
        RECT 4.000 292.080 496.000 341.680 ;
        RECT 4.400 290.680 496.000 292.080 ;
        RECT 4.000 281.200 496.000 290.680 ;
        RECT 4.000 279.800 495.600 281.200 ;
        RECT 4.000 219.320 496.000 279.800 ;
        RECT 4.000 217.920 495.600 219.320 ;
        RECT 4.000 209.120 496.000 217.920 ;
        RECT 4.400 207.720 496.000 209.120 ;
        RECT 4.000 157.440 496.000 207.720 ;
        RECT 4.000 156.040 495.600 157.440 ;
        RECT 4.000 126.160 496.000 156.040 ;
        RECT 4.400 124.760 496.000 126.160 ;
        RECT 4.000 95.560 496.000 124.760 ;
        RECT 4.000 94.160 495.600 95.560 ;
        RECT 4.000 43.200 496.000 94.160 ;
        RECT 4.400 41.800 496.000 43.200 ;
        RECT 4.000 33.680 496.000 41.800 ;
        RECT 4.000 32.280 495.600 33.680 ;
        RECT 4.000 10.715 496.000 32.280 ;
  END
END cla
END LIBRARY

