magic
tech sky130A
magscale 1 2
timestamp 1672409530
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 1104 2128 98808 97424
<< obsm2 >>
rect 1674 2139 98330 97413
<< metal3 >>
rect 0 92760 800 92880
rect 99200 87184 100000 87304
rect 0 78480 800 78600
rect 0 64200 800 64320
rect 99200 62296 100000 62416
rect 0 49920 800 50040
rect 99200 37408 100000 37528
rect 0 35640 800 35760
rect 0 21360 800 21480
rect 99200 12520 100000 12640
rect 0 7080 800 7200
<< obsm3 >>
rect 800 92960 99200 97409
rect 880 92680 99200 92960
rect 800 87384 99200 92680
rect 800 87104 99120 87384
rect 800 78680 99200 87104
rect 880 78400 99200 78680
rect 800 64400 99200 78400
rect 880 64120 99200 64400
rect 800 62496 99200 64120
rect 800 62216 99120 62496
rect 800 50120 99200 62216
rect 880 49840 99200 50120
rect 800 37608 99200 49840
rect 800 37328 99120 37608
rect 800 35840 99200 37328
rect 880 35560 99200 35840
rect 800 21560 99200 35560
rect 880 21280 99200 21560
rect 800 12720 99200 21280
rect 800 12440 99120 12720
rect 800 7280 99200 12440
rect 880 7000 99200 7280
rect 800 2143 99200 7000
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< labels >>
rlabel metal3 s 0 7080 800 7200 6 a
port 1 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 b
port 2 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 c
port 3 nsew signal output
rlabel metal3 s 0 49920 800 50040 6 d
port 4 nsew signal output
rlabel metal3 s 0 64200 800 64320 6 e
port 5 nsew signal output
rlabel metal3 s 0 78480 800 78600 6 f
port 6 nsew signal output
rlabel metal3 s 0 92760 800 92880 6 g
port 7 nsew signal output
rlabel metal3 s 99200 12520 100000 12640 6 i[0]
port 8 nsew signal input
rlabel metal3 s 99200 37408 100000 37528 6 i[1]
port 9 nsew signal input
rlabel metal3 s 99200 62296 100000 62416 6 i[2]
port 10 nsew signal input
rlabel metal3 s 99200 87184 100000 87304 6 i[3]
port 11 nsew signal input
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 12 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 13 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 13 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2648688
string GDS_FILE /home/spice/mpw8/openlane/SEVEN_SEG_DECODER/runs/22_12_30_19_37/results/signoff/SEVEN_SEG_DECODER.magic.gds
string GDS_START 117568
<< end >>

