VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO SEVEN_SEG_DECODER
  CLASS BLOCK ;
  FOREIGN SEVEN_SEG_DECODER ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN a
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END a
  PIN b
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END b
  PIN c
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END c
  PIN d
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END d
  PIN e
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END e
  PIN f
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.400 4.000 393.000 ;
    END
  END f
  PIN g
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END g
  PIN i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 62.600 500.000 63.200 ;
    END
  END i[0]
  PIN i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 187.040 500.000 187.640 ;
    END
  END i[1]
  PIN i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 311.480 500.000 312.080 ;
    END
  END i[2]
  PIN i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 435.920 500.000 436.520 ;
    END
  END i[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 5.520 10.640 494.040 487.120 ;
      LAYER met2 ;
        RECT 8.370 10.695 491.650 487.065 ;
      LAYER met3 ;
        RECT 4.000 464.800 496.000 487.045 ;
        RECT 4.400 463.400 496.000 464.800 ;
        RECT 4.000 436.920 496.000 463.400 ;
        RECT 4.000 435.520 495.600 436.920 ;
        RECT 4.000 393.400 496.000 435.520 ;
        RECT 4.400 392.000 496.000 393.400 ;
        RECT 4.000 322.000 496.000 392.000 ;
        RECT 4.400 320.600 496.000 322.000 ;
        RECT 4.000 312.480 496.000 320.600 ;
        RECT 4.000 311.080 495.600 312.480 ;
        RECT 4.000 250.600 496.000 311.080 ;
        RECT 4.400 249.200 496.000 250.600 ;
        RECT 4.000 188.040 496.000 249.200 ;
        RECT 4.000 186.640 495.600 188.040 ;
        RECT 4.000 179.200 496.000 186.640 ;
        RECT 4.400 177.800 496.000 179.200 ;
        RECT 4.000 107.800 496.000 177.800 ;
        RECT 4.400 106.400 496.000 107.800 ;
        RECT 4.000 63.600 496.000 106.400 ;
        RECT 4.000 62.200 495.600 63.600 ;
        RECT 4.000 36.400 496.000 62.200 ;
        RECT 4.400 35.000 496.000 36.400 ;
        RECT 4.000 10.715 496.000 35.000 ;
  END
END SEVEN_SEG_DECODER
END LIBRARY

