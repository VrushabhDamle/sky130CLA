magic
tech sky130A
magscale 1 2
timestamp 1672415530
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 1104 2128 98808 97424
<< obsm2 >>
rect 1582 2139 98512 97413
<< metal3 >>
rect 99200 93168 100000 93288
rect 0 91400 800 91520
rect 99200 80792 100000 80912
rect 0 74808 800 74928
rect 99200 68416 100000 68536
rect 0 58216 800 58336
rect 99200 56040 100000 56160
rect 99200 43664 100000 43784
rect 0 41624 800 41744
rect 99200 31288 100000 31408
rect 0 25032 800 25152
rect 99200 18912 100000 19032
rect 0 8440 800 8560
rect 99200 6536 100000 6656
<< obsm3 >>
rect 800 93368 99200 97409
rect 800 93088 99120 93368
rect 800 91600 99200 93088
rect 880 91320 99200 91600
rect 800 80992 99200 91320
rect 800 80712 99120 80992
rect 800 75008 99200 80712
rect 880 74728 99200 75008
rect 800 68616 99200 74728
rect 800 68336 99120 68616
rect 800 58416 99200 68336
rect 880 58136 99200 58416
rect 800 56240 99200 58136
rect 800 55960 99120 56240
rect 800 43864 99200 55960
rect 800 43584 99120 43864
rect 800 41824 99200 43584
rect 880 41544 99200 41824
rect 800 31488 99200 41544
rect 800 31208 99120 31488
rect 800 25232 99200 31208
rect 880 24952 99200 25232
rect 800 19112 99200 24952
rect 800 18832 99120 19112
rect 800 8640 99200 18832
rect 880 8360 99200 8640
rect 800 6736 99200 8360
rect 800 6456 99120 6736
rect 800 2143 99200 6456
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< labels >>
rlabel metal3 s 99200 6536 100000 6656 6 A[0]
port 1 nsew signal input
rlabel metal3 s 99200 18912 100000 19032 6 A[1]
port 2 nsew signal input
rlabel metal3 s 99200 31288 100000 31408 6 A[2]
port 3 nsew signal input
rlabel metal3 s 99200 43664 100000 43784 6 A[3]
port 4 nsew signal input
rlabel metal3 s 99200 56040 100000 56160 6 B[0]
port 5 nsew signal input
rlabel metal3 s 99200 68416 100000 68536 6 B[1]
port 6 nsew signal input
rlabel metal3 s 99200 80792 100000 80912 6 B[2]
port 7 nsew signal input
rlabel metal3 s 99200 93168 100000 93288 6 B[3]
port 8 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 S[0]
port 9 nsew signal output
rlabel metal3 s 0 25032 800 25152 6 S[1]
port 10 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 S[2]
port 11 nsew signal output
rlabel metal3 s 0 58216 800 58336 6 S[3]
port 12 nsew signal output
rlabel metal3 s 0 91400 800 91520 6 cin
port 13 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 cout
port 14 nsew signal output
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 16 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 16 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 16 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2681560
string GDS_FILE /home/spice/mpw8/openlane/cla/runs/22_12_30_21_16/results/signoff/cla.magic.gds
string GDS_START 132688
<< end >>

